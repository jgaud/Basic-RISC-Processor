library verilog;
use verilog.vl_types.all;
entity shiftLeft2_vlg_vec_tst is
end shiftLeft2_vlg_vec_tst;
