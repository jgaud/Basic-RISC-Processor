library verilog;
use verilog.vl_types.all;
entity AdderNBits_vlg_vec_tst is
end AdderNBits_vlg_vec_tst;
