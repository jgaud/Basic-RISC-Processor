library verilog;
use verilog.vl_types.all;
entity PCPlusFour_vlg_vec_tst is
end PCPlusFour_vlg_vec_tst;
